module ARM (clk, rst);
input clk;
input rst;




endmodule 